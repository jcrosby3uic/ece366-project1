module inverter(
	input A,
  	output Inv
);
	assign Inv = !A;
endmodule
